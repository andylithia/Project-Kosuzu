** sch_path:
*+ /home/andylithia/github/Project-Kosuzu/SKY130/xschem/cmos_vref/Y.Ji_JSSC2019/s2_ztat1.sch
**.subckt s2_ztat1
XQ1 GND GND v3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=5
V1 net4 GND 3
.save i(v1)
XM3 v1 v0 v0 v0 sky130_fd_pr__pfet_01v8 L=L1 W=W1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=N1 m=N1
XM1 v3 v3 net1 v2 sky130_fd_pr__pfet_01v8 L=L2 W=W2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=N2 m=N2
XM4 net1 v3 v2 v2 sky130_fd_pr__pfet_01v8 L=L2 W=W2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=N2 m=N2
XM2 v2 v2 net2 v1 sky130_fd_pr__pfet_01v8 L=L2 W=W2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=N2 m=N2
XM5 net2 v2 v1 v1 sky130_fd_pr__pfet_01v8 L=L2 W=W2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=N2 m=N2
XM6 net3 v1 v0 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 v1 net3 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.save all
.options savecurrents

.param L1=1
.param W1=20
.param N1=18

.param L2=0.5
.param W2=1
.param N2=20

.dc TEMP -20 100 1
.control
run
display
plot v0 v1 v2 v3
plot i(v1)
.endc




*.param L1=0.5
*.param W1=20
*.param N1=1
*.param L2=30
*.param W2=0.5
*.param N2=1



**** end user architecture code
**.ends
.GLOBAL GND
.end
